module ALUControl (
    input   [2:0]   ALUOp,
    input   [2:0]   funct3,
    input           funct75,
    input           OPCode5,
    output  [3:0]   ALUControlOut
);


    
endmodule