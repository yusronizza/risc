module multiplier (
    input [31:0] A,
    input [31:0] B,
    output [63:0] out
);



endmodule