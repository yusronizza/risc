module mux2x1(
    input           sel,
    input   [31:0]  inA,
    input   [31:0]  inB,
    output  [31:0]  out
);

endmodule